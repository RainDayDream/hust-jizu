/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : MAZEMAP                                                      **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module MAZEMAP( Addr,
                CLK,
                Data,
                RST,
                WE,
                R1,
                R10,
                R11,
                R12,
                R13,
                R14,
                R15,
                R16,
                R17,
                R18,
                R19,
                R2,
                R20,
                R21,
                R22,
                R23,
                R24,
                R25,
                R26,
                R27,
                R28,
                R29,
                R3,
                R30,
                R31,
                R32,
                R4,
                R5,
                R6,
                R7,
                R8,
                R9);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input[9:0]  Addr;
   input  CLK;
   input[31:0]  Data;
   input  RST;
   input  WE;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] R1;
   output[31:0] R10;
   output[31:0] R11;
   output[31:0] R12;
   output[31:0] R13;
   output[31:0] R14;
   output[31:0] R15;
   output[31:0] R16;
   output[31:0] R17;
   output[31:0] R18;
   output[31:0] R19;
   output[31:0] R2;
   output[31:0] R20;
   output[31:0] R21;
   output[31:0] R22;
   output[31:0] R23;
   output[31:0] R24;
   output[31:0] R25;
   output[31:0] R26;
   output[31:0] R27;
   output[31:0] R28;
   output[31:0] R29;
   output[31:0] R3;
   output[31:0] R30;
   output[31:0] R31;
   output[31:0] R32;
   output[31:0] R4;
   output[31:0] R5;
   output[31:0] R6;
   output[31:0] R7;
   output[31:0] R8;
   output[31:0] R9;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire[31:0] s_LOGISIM_BUS_100;
   wire[31:0] s_LOGISIM_BUS_101;
   wire[31:0] s_LOGISIM_BUS_12;
   wire[31:0] s_LOGISIM_BUS_16;
   wire[31:0] s_LOGISIM_BUS_17;
   wire[31:0] s_LOGISIM_BUS_18;
   wire[31:0] s_LOGISIM_BUS_21;
   wire[31:0] s_LOGISIM_BUS_22;
   wire[31:0] s_LOGISIM_BUS_26;
   wire[31:0] s_LOGISIM_BUS_27;
   wire[31:0] s_LOGISIM_BUS_33;
   wire[31:0] s_LOGISIM_BUS_34;
   wire[31:0] s_LOGISIM_BUS_39;
   wire[31:0] s_LOGISIM_BUS_41;
   wire[31:0] s_LOGISIM_BUS_42;
   wire[31:0] s_LOGISIM_BUS_48;
   wire[31:0] s_LOGISIM_BUS_5;
   wire[31:0] s_LOGISIM_BUS_56;
   wire[31:0] s_LOGISIM_BUS_57;
   wire[31:0] s_LOGISIM_BUS_6;
   wire[31:0] s_LOGISIM_BUS_62;
   wire[31:0] s_LOGISIM_BUS_63;
   wire[31:0] s_LOGISIM_BUS_71;
   wire[31:0] s_LOGISIM_BUS_74;
   wire[31:0] s_LOGISIM_BUS_79;
   wire[31:0] s_LOGISIM_BUS_8;
   wire[31:0] s_LOGISIM_BUS_80;
   wire[31:0] s_LOGISIM_BUS_84;
   wire[31:0] s_LOGISIM_BUS_85;
   wire[31:0] s_LOGISIM_BUS_9;
   wire[31:0] s_LOGISIM_BUS_92;
   wire[31:0] s_LOGISIM_BUS_93;
   wire[31:0] s_LOGISIM_BUS_94;
   wire[9:0] s_LOGISIM_BUS_95;
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_10;
   wire s_LOGISIM_NET_102;
   wire s_LOGISIM_NET_103;
   wire s_LOGISIM_NET_11;
   wire s_LOGISIM_NET_13;
   wire s_LOGISIM_NET_14;
   wire s_LOGISIM_NET_15;
   wire s_LOGISIM_NET_19;
   wire s_LOGISIM_NET_2;
   wire s_LOGISIM_NET_20;
   wire s_LOGISIM_NET_23;
   wire s_LOGISIM_NET_24;
   wire s_LOGISIM_NET_25;
   wire s_LOGISIM_NET_28;
   wire s_LOGISIM_NET_29;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_30;
   wire s_LOGISIM_NET_31;
   wire s_LOGISIM_NET_32;
   wire s_LOGISIM_NET_35;
   wire s_LOGISIM_NET_36;
   wire s_LOGISIM_NET_37;
   wire s_LOGISIM_NET_38;
   wire s_LOGISIM_NET_4;
   wire s_LOGISIM_NET_40;
   wire s_LOGISIM_NET_43;
   wire s_LOGISIM_NET_44;
   wire s_LOGISIM_NET_45;
   wire s_LOGISIM_NET_46;
   wire s_LOGISIM_NET_47;
   wire s_LOGISIM_NET_49;
   wire s_LOGISIM_NET_50;
   wire s_LOGISIM_NET_51;
   wire s_LOGISIM_NET_53;
   wire s_LOGISIM_NET_54;
   wire s_LOGISIM_NET_55;
   wire s_LOGISIM_NET_58;
   wire s_LOGISIM_NET_59;
   wire s_LOGISIM_NET_60;
   wire s_LOGISIM_NET_61;
   wire s_LOGISIM_NET_64;
   wire s_LOGISIM_NET_65;
   wire s_LOGISIM_NET_66;
   wire s_LOGISIM_NET_67;
   wire s_LOGISIM_NET_68;
   wire s_LOGISIM_NET_69;
   wire s_LOGISIM_NET_7;
   wire s_LOGISIM_NET_70;
   wire s_LOGISIM_NET_72;
   wire s_LOGISIM_NET_73;
   wire s_LOGISIM_NET_75;
   wire s_LOGISIM_NET_76;
   wire s_LOGISIM_NET_77;
   wire s_LOGISIM_NET_78;
   wire s_LOGISIM_NET_81;
   wire s_LOGISIM_NET_82;
   wire s_LOGISIM_NET_83;
   wire s_LOGISIM_NET_86;
   wire s_LOGISIM_NET_87;
   wire s_LOGISIM_NET_88;
   wire s_LOGISIM_NET_89;
   wire s_LOGISIM_NET_90;
   wire s_LOGISIM_NET_91;
   wire s_LOGISIM_NET_96;
   wire s_LOGISIM_NET_97;
   wire s_LOGISIM_NET_98;
   wire s_LOGISIM_NET_99;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_BUS_101[31:0]            = Data;
   assign s_LOGISIM_NET_2                    = WE;
   assign s_LOGISIM_NET_1                    = RST;
   assign s_LOGISIM_BUS_95[9:0]              = Addr;
   assign s_LOGISIM_NET_3                    = CLK;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign R23                                = s_LOGISIM_BUS_8[31:0];
   assign R5                                 = s_LOGISIM_BUS_100[31:0];
   assign R18                                = s_LOGISIM_BUS_6[31:0];
   assign R15                                = s_LOGISIM_BUS_93[31:0];
   assign R13                                = s_LOGISIM_BUS_5[31:0];
   assign R28                                = s_LOGISIM_BUS_42[31:0];
   assign R24                                = s_LOGISIM_BUS_92[31:0];
   assign R19                                = s_LOGISIM_BUS_85[31:0];
   assign R2                                 = s_LOGISIM_BUS_48[31:0];
   assign R4                                 = s_LOGISIM_BUS_12[31:0];
   assign R25                                = s_LOGISIM_BUS_17[31:0];
   assign R10                                = s_LOGISIM_BUS_57[31:0];
   assign R31                                = s_LOGISIM_BUS_94[31:0];
   assign R30                                = s_LOGISIM_BUS_9[31:0];
   assign R29                                = s_LOGISIM_BUS_22[31:0];
   assign R9                                 = s_LOGISIM_BUS_80[31:0];
   assign R3                                 = s_LOGISIM_BUS_27[31:0];
   assign R22                                = s_LOGISIM_BUS_21[31:0];
   assign R7                                 = s_LOGISIM_BUS_56[31:0];
   assign R8                                 = s_LOGISIM_BUS_33[31:0];
   assign R32                                = s_LOGISIM_BUS_74[31:0];
   assign R27                                = s_LOGISIM_BUS_63[31:0];
   assign R6                                 = s_LOGISIM_BUS_79[31:0];
   assign R16                                = s_LOGISIM_BUS_39[31:0];
   assign R11                                = s_LOGISIM_BUS_34[31:0];
   assign R12                                = s_LOGISIM_BUS_16[31:0];
   assign R26                                = s_LOGISIM_BUS_26[31:0];
   assign R1                                 = s_LOGISIM_BUS_71[31:0];
   assign R20                                = s_LOGISIM_BUS_62[31:0];
   assign R21                                = s_LOGISIM_BUS_41[31:0];
   assign R14                                = s_LOGISIM_BUS_84[31:0];
   assign R17                                = s_LOGISIM_BUS_18[31:0];

   /***************************************************************************
    ** Here all in-lined components are defined                              **
    ***************************************************************************/
   assign s_LOGISIM_NET_0 = 1'd0;

   assign s_LOGISIM_NET_61 = 1'd1;


   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   AND_GATE #(.BubblesMask(0))
      GATE_1 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_72),
              .Result(s_LOGISIM_NET_37));

   AND_GATE #(.BubblesMask(0))
      GATE_2 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_38),
              .Result(s_LOGISIM_NET_51));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_1 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_24),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_63[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   Demultiplexer_32      DEMUX_1 (.DemuxIn(s_LOGISIM_NET_61),
                                  .DemuxOut_0(s_LOGISIM_NET_40),
                                  .DemuxOut_1(s_LOGISIM_NET_38),
                                  .DemuxOut_10(s_LOGISIM_NET_72),
                                  .DemuxOut_11(s_LOGISIM_NET_54),
                                  .DemuxOut_12(s_LOGISIM_NET_28),
                                  .DemuxOut_13(s_LOGISIM_NET_35),
                                  .DemuxOut_14(s_LOGISIM_NET_102),
                                  .DemuxOut_15(s_LOGISIM_NET_90),
                                  .DemuxOut_16(s_LOGISIM_NET_91),
                                  .DemuxOut_17(s_LOGISIM_NET_73),
                                  .DemuxOut_18(s_LOGISIM_NET_49),
                                  .DemuxOut_19(s_LOGISIM_NET_29),
                                  .DemuxOut_2(s_LOGISIM_NET_86),
                                  .DemuxOut_20(s_LOGISIM_NET_13),
                                  .DemuxOut_21(s_LOGISIM_NET_103),
                                  .DemuxOut_22(s_LOGISIM_NET_81),
                                  .DemuxOut_23(s_LOGISIM_NET_58),
                                  .DemuxOut_24(s_LOGISIM_NET_64),
                                  .DemuxOut_25(s_LOGISIM_NET_43),
                                  .DemuxOut_26(s_LOGISIM_NET_23),
                                  .DemuxOut_27(s_LOGISIM_NET_15),
                                  .DemuxOut_28(s_LOGISIM_NET_96),
                                  .DemuxOut_29(s_LOGISIM_NET_75),
                                  .DemuxOut_3(s_LOGISIM_NET_67),
                                  .DemuxOut_30(s_LOGISIM_NET_50),
                                  .DemuxOut_31(s_LOGISIM_NET_30),
                                  .DemuxOut_4(s_LOGISIM_NET_44),
                                  .DemuxOut_5(s_LOGISIM_NET_65),
                                  .DemuxOut_6(s_LOGISIM_NET_20),
                                  .DemuxOut_7(s_LOGISIM_NET_97),
                                  .DemuxOut_8(s_LOGISIM_NET_66),
                                  .DemuxOut_9(s_LOGISIM_NET_89),
                                  .Enable(1'b1),
                                  .Sel(s_LOGISIM_BUS_95[4:0]));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_2 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_60),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_57[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_3 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_14),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_12[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_4 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_19),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_16[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_3 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_65),
              .Result(s_LOGISIM_NET_82));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_5 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_45),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_39[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_4 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_20),
              .Result(s_LOGISIM_NET_59));

   AND_GATE #(.BubblesMask(0))
      GATE_5 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_54),
              .Result(s_LOGISIM_NET_19));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_6 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_51),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_48[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_6 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_15),
              .Result(s_LOGISIM_NET_10));

   AND_GATE #(.BubblesMask(0))
      GATE_7 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_43),
              .Result(s_LOGISIM_NET_46));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_7 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_82),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_79[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_8 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_102),
              .Result(s_LOGISIM_NET_68));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_8 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_99),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_21[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_9 (.Input_1(s_LOGISIM_NET_2),
              .Input_2(s_LOGISIM_NET_89),
              .Result(s_LOGISIM_NET_60));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_9 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_10),
                       .D(s_LOGISIM_BUS_101[31:0]),
                       .Q(s_LOGISIM_BUS_42[31:0]),
                       .Reset(s_LOGISIM_NET_1),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_0),
                       .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_10 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_49),
               .Result(s_LOGISIM_NET_47));

   AND_GATE #(.BubblesMask(0))
      GATE_11 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_81),
               .Result(s_LOGISIM_NET_78));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_10 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_87),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_84[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_12 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_91),
               .Result(s_LOGISIM_NET_88));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_11 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_78),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_8[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_13 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_75),
               .Result(s_LOGISIM_NET_77));

   AND_GATE #(.BubblesMask(0))
      GATE_14 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_86),
               .Result(s_LOGISIM_NET_31));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_12 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_32),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_74[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_13 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_53),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_94[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_15 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_29),
               .Result(s_LOGISIM_NET_25));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_14 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_46),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_26[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_16 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_73),
               .Result(s_LOGISIM_NET_70));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_15 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_11),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_41[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_17 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_13),
               .Result(s_LOGISIM_NET_11));

   AND_GATE #(.BubblesMask(0))
      GATE_18 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_66),
               .Result(s_LOGISIM_NET_83));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_16 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_77),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_9[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_17 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_25),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_62[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_19 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_103),
               .Result(s_LOGISIM_NET_99));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_18 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_100[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_20 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_30),
               .Result(s_LOGISIM_NET_32));

   AND_GATE #(.BubblesMask(0))
      GATE_21 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_50),
               .Result(s_LOGISIM_NET_53));

   AND_GATE #(.BubblesMask(0))
      GATE_22 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_90),
               .Result(s_LOGISIM_NET_45));

   AND_GATE #(.BubblesMask(0))
      GATE_23 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_40),
               .Result(s_LOGISIM_NET_76));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_19 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_68),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_93[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_20 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_7),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_5[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_24 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_58),
               .Result(s_LOGISIM_NET_55));

   AND_GATE #(.BubblesMask(0))
      GATE_25 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_96),
               .Result(s_LOGISIM_NET_98));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_21 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_98),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_22[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_22 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_36),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_33[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_23 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_55),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_92[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_26 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_23),
               .Result(s_LOGISIM_NET_24));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_24 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_47),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_85[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_27 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_67),
               .Result(s_LOGISIM_NET_14));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_25 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_69),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_17[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_26 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_83),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_80[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_28 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_35),
               .Result(s_LOGISIM_NET_87));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_27 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_59),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_56[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_28 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_88),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_18[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_29 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_44),
               .Result(s_LOGISIM_NET_4));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_29 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_76),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_71[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_30 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_28),
               .Result(s_LOGISIM_NET_7));

   AND_GATE #(.BubblesMask(0))
      GATE_31 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_97),
               .Result(s_LOGISIM_NET_36));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_30 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_70),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_6[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_31 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_37),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_34[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_32 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_31),
                        .D(s_LOGISIM_BUS_101[31:0]),
                        .Q(s_LOGISIM_BUS_27[31:0]),
                        .Reset(s_LOGISIM_NET_1),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_0),
                        .pre(s_LOGISIM_NET_0));

   AND_GATE #(.BubblesMask(0))
      GATE_32 (.Input_1(s_LOGISIM_NET_2),
               .Input_2(s_LOGISIM_NET_64),
               .Result(s_LOGISIM_NET_69));



endmodule
