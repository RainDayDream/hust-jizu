/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : ROM_IRPLACE                                                  **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module ROM_IRPLACE( Address,
                    Data);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input[9:0]  Address;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] Data;
   reg[31:0] Data;

   always @ (Address)
   begin
      case(Address)
         0 : Data = 1258291311;
         1 : Data = 403249251;
         2 : Data = 268960567;
         3 : Data = 1245971;
         4 : Data = 6299683;
         5 : Data = 268960567;
         6 : Data = 197395;
         7 : Data = 6300195;
         8 : Data = 520651575;
         9 : Data = -470613229;
         10 : Data = 6300707;
         11 : Data = 17302327;
         12 : Data = 537068307;
         13 : Data = 6301219;
         14 : Data = -519568585;
         15 : Data = 537068307;
         16 : Data = 6301731;
         17 : Data = 16810807;
         18 : Data = -8191213;
         19 : Data = 6302243;
         20 : Data = 16794423;
         21 : Data = 197395;
         22 : Data = 6302755;
         23 : Data = -16760009;
         24 : Data = 197395;
         25 : Data = 6303267;
         26 : Data = 269472567;
         27 : Data = -8191213;
         28 : Data = 39854115;
         29 : Data = 268964663;
         30 : Data = -2147286253;
         31 : Data = 39854627;
         32 : Data = 268964663;
         33 : Data = -2147286253;
         34 : Data = 39855139;
         35 : Data = 335024951;
         36 : Data = -2147286253;
         37 : Data = 39855651;
         38 : Data = 302777143;
         39 : Data = -1879899373;
         40 : Data = 39856163;
         41 : Data = 302646071;
         42 : Data = 134415123;
         43 : Data = 39856675;
         44 : Data = 305791799;
         45 : Data = 134415123;
         46 : Data = 39857187;
         47 : Data = 270664503;
         48 : Data = 134415123;
         49 : Data = 39857699;
         50 : Data = 270730039;
         51 : Data = -268238061;
         52 : Data = 73408547;
         53 : Data = 300024631;
         54 : Data = 8586003;
         55 : Data = 73409059;
         56 : Data = 285213495;
         57 : Data = 8586003;
         58 : Data = 73409571;
         59 : Data = 285213495;
         60 : Data = 8586003;
         61 : Data = 73410083;
         62 : Data = -12586185;
         63 : Data = 2139292435;
         64 : Data = 73410595;
         65 : Data = 18879287;
         66 : Data = -2147286253;
         67 : Data = 73411107;
         68 : Data = 18879287;
         69 : Data = -2147286253;
         70 : Data = 73411619;
         71 : Data = 18879287;
         72 : Data = -2147286253;
         73 : Data = 73412131;
         74 : Data = -114425033;
         75 : Data = 1072890643;
         76 : Data = 106962979;
         77 : Data = 1091048247;
         78 : Data = -2147286253;
         79 : Data = 106963491;
         80 : Data = 1091048247;
         81 : Data = -2147286253;
         82 : Data = 106964003;
         83 : Data = 1091048247;
         84 : Data = -2147286253;
         85 : Data = 106964515;
         86 : Data = 536363831;
         87 : Data = -259849453;
         88 : Data = 106965027;
         89 : Data = 9015;
         90 : Data = 8586003;
         91 : Data = 106965539;
         92 : Data = 9015;
         93 : Data = 8586003;
         94 : Data = 106966051;
         95 : Data = 536806199;
         96 : Data = 8586003;
         97 : Data = 106966563;
         98 : Data = 35653779;
         99 : Data = 115;
         100 : Data = 1050899;
         101 : Data = 2097267;
         102 : Data = 403249251;
         103 : Data = 383845175;
         104 : Data = -7142637;
         105 : Data = 6299683;
         106 : Data = 268702519;
         107 : Data = -528284909;
         108 : Data = 6300195;
         109 : Data = 268903223;
         110 : Data = 69403411;
         111 : Data = 6300707;
         112 : Data = 284967735;
         113 : Data = -8191213;
         114 : Data = 6301219;
         115 : Data = 1200951;
         116 : Data = 153289491;
         117 : Data = 6301731;
         118 : Data = -15428809;
         119 : Data = 178455315;
         120 : Data = 6302243;
         121 : Data = 5919543;
         122 : Data = 207815443;
         123 : Data = 6302755;
         124 : Data = -2854089;
         125 : Data = 1240662803;
         126 : Data = 6303267;
         127 : Data = 135283511;
         128 : Data = 1252197139;
         129 : Data = 39854115;
         130 : Data = 1511564087;
         131 : Data = 1834156819;
         132 : Data = 39854627;
         133 : Data = -1525415113;
         134 : Data = 1252197139;
         135 : Data = 39855139;
         136 : Data = 1610613559;
         137 : Data = -806157549;
         138 : Data = 39855651;
         139 : Data = 277394231;
         140 : Data = 177406739;
         141 : Data = 39856163;
         142 : Data = 341119799;
         143 : Data = 142803731;
         144 : Data = 39856675;
         145 : Data = -199081161;
         146 : Data = 1956840211;
         147 : Data = 39857187;
         148 : Data = 100623159;
         149 : Data = 1117979411;
         150 : Data = 39857699;
         151 : Data = -8109257;
         152 : Data = 1352860435;
         153 : Data = 73408547;
         154 : Data = 289891127;
         155 : Data = -728562925;
         156 : Data = 73409059;
         157 : Data = 1226855223;
         158 : Data = 617808659;
         159 : Data = 73409571;
         160 : Data = -14691529;
         161 : Data = 347276051;
         162 : Data = 73410083;
         163 : Data = 542122807;
         164 : Data = -40697069;
         165 : Data = 73410595;
         166 : Data = 278225719;
         167 : Data = -1986854125;
         168 : Data = 73411107;
         169 : Data = -921423049;
         170 : Data = 1389560595;
         171 : Data = 73411619;
         172 : Data = 536081207;
         173 : Data = 546505491;
         174 : Data = 73412131;
         175 : Data = -2146229449;
         176 : Data = 1609761555;
         177 : Data = 106962979;
         178 : Data = -2138668233;
         179 : Data = 1212351251;
         180 : Data = 106963491;
         181 : Data = -1610722505;
         182 : Data = 1279460115;
         183 : Data = 106964003;
         184 : Data = 4207415;
         185 : Data = 1551041299;
         186 : Data = 106964515;
         187 : Data = 809784119;
         188 : Data = 690160403;
         189 : Data = 106965027;
         190 : Data = -58813641;
         191 : Data = 1607664403;
         192 : Data = 106965539;
         193 : Data = 1276257079;
         194 : Data = -2002582765;
         195 : Data = 106966051;
         196 : Data = 54071;
         197 : Data = 75694867;
         198 : Data = 106966563;
         199 : Data = 35653779;
         200 : Data = 115;
         201 : Data = 1050899;
         202 : Data = 2097267;
         203 : Data = 67701347;
         204 : Data = 32506643;
         205 : Data = 375654499;
         206 : Data = 1049363;
         207 : Data = 6554547;
         208 : Data = 7544371;
         209 : Data = 2399891;
         210 : Data = 962307;
         211 : Data = 30375859;
         212 : Data = 336566883;
         213 : Data = 6554675;
         214 : Data = 30371635;
         215 : Data = 1990163;
         216 : Data = 30363443;
         217 : Data = 32415779;
         218 : Data = 35653779;
         219 : Data = 115;
         220 : Data = 32506771;
         221 : Data = 7603299;
         222 : Data = 2097267;
         223 : Data = 544508003;
         224 : Data = 2097267;
         225 : Data = 67701347;
         226 : Data = 915;
         227 : Data = 276040803;
         228 : Data = 1049363;
         229 : Data = 1080296371;
         230 : Data = 7544371;
         231 : Data = 2399891;
         232 : Data = 962307;
         233 : Data = 30375859;
         234 : Data = 235904611;
         235 : Data = 1080296499;
         236 : Data = 30371635;
         237 : Data = 1973779;
         238 : Data = 30363443;
         239 : Data = 32415779;
         240 : Data = 35653779;
         241 : Data = 115;
         242 : Data = 32506771;
         243 : Data = 7603299;
         244 : Data = 2097267;
         245 : Data = 443845731;
         246 : Data = 2097267;
         247 : Data = 101253219;
         248 : Data = 32506771;
         249 : Data = 208961635;
         250 : Data = 1049363;
         251 : Data = 8592947;
         252 : Data = 6587315;
         253 : Data = 2334355;
         254 : Data = 962307;
         255 : Data = 30375859;
         256 : Data = 168792675;
         257 : Data = 6587571;
         258 : Data = 30371635;
         259 : Data = 32415779;
         260 : Data = 4195219;
         261 : Data = 1082035891;
         262 : Data = 962307;
         263 : Data = 30363443;
         264 : Data = 32415779;
         265 : Data = 35653779;
         266 : Data = 115;
         267 : Data = 32506771;
         268 : Data = 7603299;
         269 : Data = 2097267;
         270 : Data = 343181923;
         271 : Data = 2097267;
         272 : Data = 915;
         273 : Data = 75042403;
         274 : Data = 915;
         275 : Data = 74746979;
         276 : Data = 1049363;
         277 : Data = 8592947;
         278 : Data = 1080329139;
         279 : Data = 2334355;
         280 : Data = 962307;
         281 : Data = 30375859;
         282 : Data = 34578019;
         283 : Data = 1080329395;
         284 : Data = 30371635;
         285 : Data = 32415779;
         286 : Data = 5148307;
         287 : Data = 962307;
         288 : Data = 30363443;
         289 : Data = 32415779;
         290 : Data = 35653779;
         291 : Data = 115;
         292 : Data = 32506771;
         293 : Data = 7603299;
         294 : Data = 2097267;
         295 : Data = 242518115;
         296 : Data = 2097267;
         297 : Data = 104858899;
         298 : Data = 115;
         299 : Data = 2097267;
         300 : Data = 1043;
         301 : Data = 1171;
         302 : Data = 285770551;
         303 : Data = -813497581;
         304 : Data = 6302755;
         305 : Data = 454300471;
         306 : Data = -2013068525;
         307 : Data = 6303267;
         308 : Data = 356389687;
         309 : Data = 260244243;
         310 : Data = 39854115;
         311 : Data = 287449911;
         312 : Data = 134415123;
         313 : Data = 39854627;
         314 : Data = 287474487;
         315 : Data = -813497581;
         316 : Data = 39855139;
         317 : Data = 101602103;
         318 : Data = -368901357;
         319 : Data = 39856675;
         320 : Data = 34124599;
         321 : Data = -1979514093;
         322 : Data = 39857187;
         323 : Data = 34534199;
         324 : Data = -469564653;
         325 : Data = 39857699;
         326 : Data = 34120503;
         327 : Data = 604177171;
         328 : Data = 73408547;
         329 : Data = 122598199;
         330 : Data = -469564653;
         331 : Data = 73409059;
         332 : Data = 118117175;
         333 : Data = -335346925;
         334 : Data = 73410595;
         335 : Data = 17478455;
         336 : Data = -1442643181;
         337 : Data = 73411107;
         338 : Data = 118420279;
         339 : Data = -368901357;
         340 : Data = 73411619;
         341 : Data = 67810103;
         342 : Data = -905772269;
         343 : Data = 73412131;
         344 : Data = 122336055;
         345 : Data = -1409088749;
         346 : Data = 106962979;
         347 : Data = 35653779;
         348 : Data = 115;
         349 : Data = 19;
         350 : Data = 19;
         351 : Data = 19;
         352 : Data = 19;
         353 : Data = 19;
         354 : Data = -18878353;
         355 : Data = 1051027;
         356 : Data = 787;
         357 : Data = 6299683;
         358 : Data = 787;
         359 : Data = 6300195;
         360 : Data = 787;
         361 : Data = 6300707;
         362 : Data = 787;
         363 : Data = 6301219;
         364 : Data = 787;
         365 : Data = 6301731;
         366 : Data = 787;
         367 : Data = 6302243;
         368 : Data = 787;
         369 : Data = 6302755;
         370 : Data = 787;
         371 : Data = 6303267;
         372 : Data = 787;
         373 : Data = 39854115;
         374 : Data = 787;
         375 : Data = 39854627;
         376 : Data = 787;
         377 : Data = 39855139;
         378 : Data = 787;
         379 : Data = 39855651;
         380 : Data = 787;
         381 : Data = 39856163;
         382 : Data = 1970762551;
         383 : Data = 1998783251;
         384 : Data = 39856675;
         385 : Data = 1162105655;
         386 : Data = 1143145235;
         387 : Data = 39857187;
         388 : Data = 1967420215;
         389 : Data = 1998783251;
         390 : Data = 39857699;
         391 : Data = 356795191;
         392 : Data = 285410067;
         393 : Data = 73408547;
         394 : Data = 2004316983;
         395 : Data = 1998783251;
         396 : Data = 73409059;
         397 : Data = 787;
         398 : Data = 73409571;
         399 : Data = 787;
         400 : Data = 73410083;
         401 : Data = 787;
         402 : Data = 73410595;
         403 : Data = 787;
         404 : Data = 73411107;
         405 : Data = 787;
         406 : Data = 73411619;
         407 : Data = 787;
         408 : Data = 73412131;
         409 : Data = 787;
         410 : Data = 106962979;
         411 : Data = 787;
         412 : Data = 106963491;
         413 : Data = 787;
         414 : Data = 106964003;
         415 : Data = 787;
         416 : Data = 106964515;
         417 : Data = 787;
         418 : Data = 106965027;
         419 : Data = 787;
         420 : Data = 106965539;
         421 : Data = 787;
         422 : Data = 106966051;
         423 : Data = 787;
         424 : Data = 106966563;
         425 : Data = 35653779;
         426 : Data = 115;
         427 : Data = -325062545;
         default : Data = 0;
      endcase
   end

endmodule
