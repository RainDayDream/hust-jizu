/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : DISPLAY                                                      **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module DISPLAY( A1,
                A10,
                A11,
                A12,
                A13,
                A14,
                A15,
                A16,
                A17,
                A18,
                A19,
                A2,
                A20,
                A21,
                A22,
                A23,
                A24,
                A25,
                A26,
                A27,
                A28,
                A29,
                A3,
                A30,
                A31,
                A32,
                A4,
                A5,
                A6,
                A7,
                A8,
                A9,
                CLK,
                RST,
                WE,
                R13,
                R1,
                R10,
                R11,
                R12,
                R14,
                R15,
                R16,
                R17,
                R18,
                R19,
                R2,
                R20,
                R21,
                R22,
                R23,
                R24,
                R25,
                R26,
                R27,
                R28,
                R29,
                R3,
                R30,
                R31,
                R32,
                R4,
                R5,
                R6,
                R7,
                R8,
                R9);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input[31:0]  A1;
   input[31:0]  A10;
   input[31:0]  A11;
   input[31:0]  A12;
   input[31:0]  A13;
   input[31:0]  A14;
   input[31:0]  A15;
   input[31:0]  A16;
   input[31:0]  A17;
   input[31:0]  A18;
   input[31:0]  A19;
   input[31:0]  A2;
   input[31:0]  A20;
   input[31:0]  A21;
   input[31:0]  A22;
   input[31:0]  A23;
   input[31:0]  A24;
   input[31:0]  A25;
   input[31:0]  A26;
   input[31:0]  A27;
   input[31:0]  A28;
   input[31:0]  A29;
   input[31:0]  A3;
   input[31:0]  A30;
   input[31:0]  A31;
   input[31:0]  A32;
   input[31:0]  A4;
   input[31:0]  A5;
   input[31:0]  A6;
   input[31:0]  A7;
   input[31:0]  A8;
   input[31:0]  A9;
   input  CLK;
   input  RST;
   input  WE;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output[31:0] R13;
   output[31:0] R1;
   output[31:0] R10;
   output[31:0] R11;
   output[31:0] R12;
   output[31:0] R14;
   output[31:0] R15;
   output[31:0] R16;
   output[31:0] R17;
   output[31:0] R18;
   output[31:0] R19;
   output[31:0] R2;
   output[31:0] R20;
   output[31:0] R21;
   output[31:0] R22;
   output[31:0] R23;
   output[31:0] R24;
   output[31:0] R25;
   output[31:0] R26;
   output[31:0] R27;
   output[31:0] R28;
   output[31:0] R29;
   output[31:0] R3;
   output[31:0] R30;
   output[31:0] R31;
   output[31:0] R32;
   output[31:0] R4;
   output[31:0] R5;
   output[31:0] R6;
   output[31:0] R7;
   output[31:0] R8;
   output[31:0] R9;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire[31:0] s_LOGISIM_BUS_0;
   wire[31:0] s_LOGISIM_BUS_10;
   wire[31:0] s_LOGISIM_BUS_11;
   wire[31:0] s_LOGISIM_BUS_12;
   wire[31:0] s_LOGISIM_BUS_13;
   wire[31:0] s_LOGISIM_BUS_14;
   wire[31:0] s_LOGISIM_BUS_15;
   wire[31:0] s_LOGISIM_BUS_16;
   wire[31:0] s_LOGISIM_BUS_17;
   wire[31:0] s_LOGISIM_BUS_18;
   wire[31:0] s_LOGISIM_BUS_19;
   wire[31:0] s_LOGISIM_BUS_2;
   wire[31:0] s_LOGISIM_BUS_20;
   wire[31:0] s_LOGISIM_BUS_21;
   wire[31:0] s_LOGISIM_BUS_22;
   wire[31:0] s_LOGISIM_BUS_23;
   wire[31:0] s_LOGISIM_BUS_24;
   wire[31:0] s_LOGISIM_BUS_25;
   wire[31:0] s_LOGISIM_BUS_26;
   wire[31:0] s_LOGISIM_BUS_27;
   wire[31:0] s_LOGISIM_BUS_28;
   wire[31:0] s_LOGISIM_BUS_29;
   wire[31:0] s_LOGISIM_BUS_30;
   wire[31:0] s_LOGISIM_BUS_31;
   wire[31:0] s_LOGISIM_BUS_32;
   wire[31:0] s_LOGISIM_BUS_33;
   wire[31:0] s_LOGISIM_BUS_34;
   wire[31:0] s_LOGISIM_BUS_35;
   wire[31:0] s_LOGISIM_BUS_36;
   wire[31:0] s_LOGISIM_BUS_37;
   wire[31:0] s_LOGISIM_BUS_38;
   wire[31:0] s_LOGISIM_BUS_39;
   wire[31:0] s_LOGISIM_BUS_40;
   wire[31:0] s_LOGISIM_BUS_41;
   wire[31:0] s_LOGISIM_BUS_42;
   wire[31:0] s_LOGISIM_BUS_43;
   wire[31:0] s_LOGISIM_BUS_44;
   wire[31:0] s_LOGISIM_BUS_45;
   wire[31:0] s_LOGISIM_BUS_46;
   wire[31:0] s_LOGISIM_BUS_47;
   wire[31:0] s_LOGISIM_BUS_48;
   wire[31:0] s_LOGISIM_BUS_49;
   wire[31:0] s_LOGISIM_BUS_5;
   wire[31:0] s_LOGISIM_BUS_50;
   wire[31:0] s_LOGISIM_BUS_51;
   wire[31:0] s_LOGISIM_BUS_52;
   wire[31:0] s_LOGISIM_BUS_53;
   wire[31:0] s_LOGISIM_BUS_54;
   wire[31:0] s_LOGISIM_BUS_55;
   wire[31:0] s_LOGISIM_BUS_56;
   wire[31:0] s_LOGISIM_BUS_57;
   wire[31:0] s_LOGISIM_BUS_58;
   wire[31:0] s_LOGISIM_BUS_59;
   wire[31:0] s_LOGISIM_BUS_60;
   wire[31:0] s_LOGISIM_BUS_61;
   wire[31:0] s_LOGISIM_BUS_62;
   wire[31:0] s_LOGISIM_BUS_63;
   wire[31:0] s_LOGISIM_BUS_64;
   wire[31:0] s_LOGISIM_BUS_65;
   wire[31:0] s_LOGISIM_BUS_66;
   wire[31:0] s_LOGISIM_BUS_67;
   wire[31:0] s_LOGISIM_BUS_7;
   wire[31:0] s_LOGISIM_BUS_8;
   wire[31:0] s_LOGISIM_BUS_9;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_4;
   wire s_LOGISIM_NET_6;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_NET_6                    = RST;
   assign s_LOGISIM_NET_4                    = WE;
   assign s_LOGISIM_BUS_44[31:0]             = A4;
   assign s_LOGISIM_BUS_50[31:0]             = A23;
   assign s_LOGISIM_BUS_8[31:0]              = A32;
   assign s_LOGISIM_BUS_54[31:0]             = A27;
   assign s_LOGISIM_BUS_41[31:0]             = A15;
   assign s_LOGISIM_BUS_13[31:0]             = A17;
   assign s_LOGISIM_BUS_31[31:0]             = A18;
   assign s_LOGISIM_BUS_11[31:0]             = A13;
   assign s_LOGISIM_BUS_64[31:0]             = A24;
   assign s_LOGISIM_BUS_56[31:0]             = A16;
   assign s_LOGISIM_BUS_0[31:0]              = A28;
   assign s_LOGISIM_BUS_23[31:0]             = A10;
   assign s_LOGISIM_NET_3                    = CLK;
   assign s_LOGISIM_BUS_35[31:0]             = A22;
   assign s_LOGISIM_BUS_63[31:0]             = A1;
   assign s_LOGISIM_BUS_18[31:0]             = A21;
   assign s_LOGISIM_BUS_19[31:0]             = A6;
   assign s_LOGISIM_BUS_58[31:0]             = A31;
   assign s_LOGISIM_BUS_29[31:0]             = A3;
   assign s_LOGISIM_BUS_67[31:0]             = A5;
   assign s_LOGISIM_BUS_60[31:0]             = A20;
   assign s_LOGISIM_BUS_39[31:0]             = A26;
   assign s_LOGISIM_BUS_22[31:0]             = A25;
   assign s_LOGISIM_BUS_33[31:0]             = A7;
   assign s_LOGISIM_BUS_7[31:0]              = A9;
   assign s_LOGISIM_BUS_52[31:0]             = A12;
   assign s_LOGISIM_BUS_26[31:0]             = A29;
   assign s_LOGISIM_BUS_48[31:0]             = A8;
   assign s_LOGISIM_BUS_37[31:0]             = A11;
   assign s_LOGISIM_BUS_46[31:0]             = A19;
   assign s_LOGISIM_BUS_43[31:0]             = A30;
   assign s_LOGISIM_BUS_27[31:0]             = A14;
   assign s_LOGISIM_BUS_15[31:0]             = A2;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign R7                                 = s_LOGISIM_BUS_49[31:0];
   assign R27                                = s_LOGISIM_BUS_2[31:0];
   assign R20                                = s_LOGISIM_BUS_12[31:0];
   assign R9                                 = s_LOGISIM_BUS_21[31:0];
   assign R30                                = s_LOGISIM_BUS_59[31:0];
   assign R2                                 = s_LOGISIM_BUS_30[31:0];
   assign R19                                = s_LOGISIM_BUS_62[31:0];
   assign R15                                = s_LOGISIM_BUS_57[31:0];
   assign R13                               = s_LOGISIM_BUS_25[31:0];
   assign R23                                = s_LOGISIM_BUS_66[31:0];
   assign R22                                = s_LOGISIM_BUS_51[31:0];
   assign R10                                = s_LOGISIM_BUS_38[31:0];
   assign R18                                = s_LOGISIM_BUS_47[31:0];
   assign R1                                 = s_LOGISIM_BUS_14[31:0];
   assign R25                                = s_LOGISIM_BUS_36[31:0];
   assign R29                                = s_LOGISIM_BUS_40[31:0];
   assign R8                                 = s_LOGISIM_BUS_65[31:0];
   assign R14                                = s_LOGISIM_BUS_42[31:0];
   assign R5                                 = s_LOGISIM_BUS_17[31:0];
   assign R28                                = s_LOGISIM_BUS_20[31:0];
   assign R24                                = s_LOGISIM_BUS_16[31:0];
   assign R11                                = s_LOGISIM_BUS_53[31:0];
   assign R3                                 = s_LOGISIM_BUS_45[31:0];
   assign R12                                = s_LOGISIM_BUS_5[31:0];
   assign R17                                = s_LOGISIM_BUS_28[31:0];
   assign R21                                = s_LOGISIM_BUS_32[31:0];
   assign R32                                = s_LOGISIM_BUS_24[31:0];
   assign R6                                 = s_LOGISIM_BUS_34[31:0];
   assign R16                                = s_LOGISIM_BUS_10[31:0];
   assign R26                                = s_LOGISIM_BUS_55[31:0];
   assign R31                                = s_LOGISIM_BUS_9[31:0];
   assign R4                                 = s_LOGISIM_BUS_61[31:0];

   /***************************************************************************
    ** Here all in-lined components are defined                              **
    ***************************************************************************/
   assign s_LOGISIM_NET_1 = 1'd0;


   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_1 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_29[31:0]),
                       .Q(s_LOGISIM_BUS_45[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_2 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_67[31:0]),
                       .Q(s_LOGISIM_BUS_17[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_3 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_0[31:0]),
                       .Q(s_LOGISIM_BUS_20[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_4 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_7[31:0]),
                       .Q(s_LOGISIM_BUS_21[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_5 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_54[31:0]),
                       .Q(s_LOGISIM_BUS_2[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_6 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_19[31:0]),
                       .Q(s_LOGISIM_BUS_34[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_7 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_27[31:0]),
                       .Q(s_LOGISIM_BUS_42[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_8 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_44[31:0]),
                       .Q(s_LOGISIM_BUS_61[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_9 (.Clock(s_LOGISIM_NET_3),
                       .ClockEnable(s_LOGISIM_NET_4),
                       .D(s_LOGISIM_BUS_13[31:0]),
                       .Q(s_LOGISIM_BUS_28[31:0]),
                       .Reset(s_LOGISIM_NET_6),
                       .Tick(1'b1),
                       .cs(s_LOGISIM_NET_1),
                       .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_10 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_11[31:0]),
                        .Q(s_LOGISIM_BUS_25[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_11 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_39[31:0]),
                        .Q(s_LOGISIM_BUS_55[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_12 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_37[31:0]),
                        .Q(s_LOGISIM_BUS_53[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_13 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_43[31:0]),
                        .Q(s_LOGISIM_BUS_59[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_14 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_48[31:0]),
                        .Q(s_LOGISIM_BUS_65[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_15 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_52[31:0]),
                        .Q(s_LOGISIM_BUS_5[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_16 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_50[31:0]),
                        .Q(s_LOGISIM_BUS_66[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_17 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_58[31:0]),
                        .Q(s_LOGISIM_BUS_9[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_18 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_26[31:0]),
                        .Q(s_LOGISIM_BUS_40[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_19 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_63[31:0]),
                        .Q(s_LOGISIM_BUS_14[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_20 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_31[31:0]),
                        .Q(s_LOGISIM_BUS_47[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_21 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_22[31:0]),
                        .Q(s_LOGISIM_BUS_36[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_22 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_64[31:0]),
                        .Q(s_LOGISIM_BUS_16[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_23 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_8[31:0]),
                        .Q(s_LOGISIM_BUS_24[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_24 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_56[31:0]),
                        .Q(s_LOGISIM_BUS_10[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_25 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_35[31:0]),
                        .Q(s_LOGISIM_BUS_51[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_26 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_60[31:0]),
                        .Q(s_LOGISIM_BUS_12[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_27 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_15[31:0]),
                        .Q(s_LOGISIM_BUS_30[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_28 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_33[31:0]),
                        .Q(s_LOGISIM_BUS_49[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_29 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_23[31:0]),
                        .Q(s_LOGISIM_BUS_38[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_30 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_46[31:0]),
                        .Q(s_LOGISIM_BUS_62[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_31 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_18[31:0]),
                        .Q(s_LOGISIM_BUS_32[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));

   REGISTER_FLIP_FLOP #(.ActiveLevel(1),
                        .NrOfBits(32))
      REGISTER_FILE_32 (.Clock(s_LOGISIM_NET_3),
                        .ClockEnable(s_LOGISIM_NET_4),
                        .D(s_LOGISIM_BUS_41[31:0]),
                        .Q(s_LOGISIM_BUS_57[31:0]),
                        .Reset(s_LOGISIM_NET_6),
                        .Tick(1'b1),
                        .cs(s_LOGISIM_NET_1),
                        .pre(s_LOGISIM_NET_1));



endmodule
