/******************************************************************************
 ** Logisim goes FPGA automatic generated Verilog code                       **
 **                                                                          **
 ** Component : CONTROLSIGNAL                                                **
 **                                                                          **
 ******************************************************************************/

`timescale 1ns/1ps
module CONTROLSIGNAL( F12,
                      F13,
                      F14,
                      F25,
                      F30,
                      OP2,
                      OP3,
                      OP4,
                      OP5,
                      OP6,
                      ALU_SRC,
                      BEQ,
                      BNE,
                      CSR,
                      JAL,
                      JALR,
                      MemToReg,
                      MemWrite,
                      RegWrite,
                      S_Type,
                      ecall,
                      half);

   /***************************************************************************
    ** Here the inputs are defined                                           **
    ***************************************************************************/
   input  F12;
   input  F13;
   input  F14;
   input  F25;
   input  F30;
   input  OP2;
   input  OP3;
   input  OP4;
   input  OP5;
   input  OP6;

   /***************************************************************************
    ** Here the outputs are defined                                          **
    ***************************************************************************/
   output ALU_SRC;
   output BEQ;
   output BNE;
   output CSR;
   output JAL;
   output JALR;
   output MemToReg;
   output MemWrite;
   output RegWrite;
   output S_Type;
   output ecall;
   output half;

   /***************************************************************************
    ** Here the internal wires are defined                                   **
    ***************************************************************************/
   wire s_LOGISIM_NET_0;
   wire s_LOGISIM_NET_1;
   wire s_LOGISIM_NET_10;
   wire s_LOGISIM_NET_100;
   wire s_LOGISIM_NET_101;
   wire s_LOGISIM_NET_102;
   wire s_LOGISIM_NET_103;
   wire s_LOGISIM_NET_104;
   wire s_LOGISIM_NET_105;
   wire s_LOGISIM_NET_106;
   wire s_LOGISIM_NET_107;
   wire s_LOGISIM_NET_108;
   wire s_LOGISIM_NET_109;
   wire s_LOGISIM_NET_11;
   wire s_LOGISIM_NET_110;
   wire s_LOGISIM_NET_111;
   wire s_LOGISIM_NET_112;
   wire s_LOGISIM_NET_113;
   wire s_LOGISIM_NET_114;
   wire s_LOGISIM_NET_115;
   wire s_LOGISIM_NET_116;
   wire s_LOGISIM_NET_117;
   wire s_LOGISIM_NET_118;
   wire s_LOGISIM_NET_119;
   wire s_LOGISIM_NET_12;
   wire s_LOGISIM_NET_120;
   wire s_LOGISIM_NET_121;
   wire s_LOGISIM_NET_122;
   wire s_LOGISIM_NET_123;
   wire s_LOGISIM_NET_124;
   wire s_LOGISIM_NET_125;
   wire s_LOGISIM_NET_126;
   wire s_LOGISIM_NET_127;
   wire s_LOGISIM_NET_128;
   wire s_LOGISIM_NET_129;
   wire s_LOGISIM_NET_13;
   wire s_LOGISIM_NET_130;
   wire s_LOGISIM_NET_131;
   wire s_LOGISIM_NET_132;
   wire s_LOGISIM_NET_133;
   wire s_LOGISIM_NET_134;
   wire s_LOGISIM_NET_135;
   wire s_LOGISIM_NET_136;
   wire s_LOGISIM_NET_137;
   wire s_LOGISIM_NET_138;
   wire s_LOGISIM_NET_139;
   wire s_LOGISIM_NET_14;
   wire s_LOGISIM_NET_140;
   wire s_LOGISIM_NET_141;
   wire s_LOGISIM_NET_142;
   wire s_LOGISIM_NET_143;
   wire s_LOGISIM_NET_144;
   wire s_LOGISIM_NET_145;
   wire s_LOGISIM_NET_146;
   wire s_LOGISIM_NET_147;
   wire s_LOGISIM_NET_148;
   wire s_LOGISIM_NET_149;
   wire s_LOGISIM_NET_15;
   wire s_LOGISIM_NET_150;
   wire s_LOGISIM_NET_151;
   wire s_LOGISIM_NET_152;
   wire s_LOGISIM_NET_153;
   wire s_LOGISIM_NET_154;
   wire s_LOGISIM_NET_155;
   wire s_LOGISIM_NET_156;
   wire s_LOGISIM_NET_157;
   wire s_LOGISIM_NET_158;
   wire s_LOGISIM_NET_159;
   wire s_LOGISIM_NET_16;
   wire s_LOGISIM_NET_160;
   wire s_LOGISIM_NET_161;
   wire s_LOGISIM_NET_162;
   wire s_LOGISIM_NET_163;
   wire s_LOGISIM_NET_164;
   wire s_LOGISIM_NET_165;
   wire s_LOGISIM_NET_166;
   wire s_LOGISIM_NET_167;
   wire s_LOGISIM_NET_168;
   wire s_LOGISIM_NET_169;
   wire s_LOGISIM_NET_17;
   wire s_LOGISIM_NET_170;
   wire s_LOGISIM_NET_171;
   wire s_LOGISIM_NET_172;
   wire s_LOGISIM_NET_173;
   wire s_LOGISIM_NET_174;
   wire s_LOGISIM_NET_175;
   wire s_LOGISIM_NET_176;
   wire s_LOGISIM_NET_177;
   wire s_LOGISIM_NET_178;
   wire s_LOGISIM_NET_179;
   wire s_LOGISIM_NET_18;
   wire s_LOGISIM_NET_180;
   wire s_LOGISIM_NET_181;
   wire s_LOGISIM_NET_182;
   wire s_LOGISIM_NET_183;
   wire s_LOGISIM_NET_184;
   wire s_LOGISIM_NET_185;
   wire s_LOGISIM_NET_186;
   wire s_LOGISIM_NET_187;
   wire s_LOGISIM_NET_188;
   wire s_LOGISIM_NET_189;
   wire s_LOGISIM_NET_19;
   wire s_LOGISIM_NET_190;
   wire s_LOGISIM_NET_191;
   wire s_LOGISIM_NET_192;
   wire s_LOGISIM_NET_193;
   wire s_LOGISIM_NET_194;
   wire s_LOGISIM_NET_195;
   wire s_LOGISIM_NET_196;
   wire s_LOGISIM_NET_197;
   wire s_LOGISIM_NET_198;
   wire s_LOGISIM_NET_199;
   wire s_LOGISIM_NET_2;
   wire s_LOGISIM_NET_20;
   wire s_LOGISIM_NET_200;
   wire s_LOGISIM_NET_201;
   wire s_LOGISIM_NET_202;
   wire s_LOGISIM_NET_203;
   wire s_LOGISIM_NET_204;
   wire s_LOGISIM_NET_205;
   wire s_LOGISIM_NET_206;
   wire s_LOGISIM_NET_207;
   wire s_LOGISIM_NET_208;
   wire s_LOGISIM_NET_209;
   wire s_LOGISIM_NET_21;
   wire s_LOGISIM_NET_210;
   wire s_LOGISIM_NET_211;
   wire s_LOGISIM_NET_212;
   wire s_LOGISIM_NET_213;
   wire s_LOGISIM_NET_214;
   wire s_LOGISIM_NET_215;
   wire s_LOGISIM_NET_216;
   wire s_LOGISIM_NET_217;
   wire s_LOGISIM_NET_218;
   wire s_LOGISIM_NET_219;
   wire s_LOGISIM_NET_22;
   wire s_LOGISIM_NET_220;
   wire s_LOGISIM_NET_221;
   wire s_LOGISIM_NET_222;
   wire s_LOGISIM_NET_223;
   wire s_LOGISIM_NET_224;
   wire s_LOGISIM_NET_225;
   wire s_LOGISIM_NET_226;
   wire s_LOGISIM_NET_227;
   wire s_LOGISIM_NET_228;
   wire s_LOGISIM_NET_229;
   wire s_LOGISIM_NET_23;
   wire s_LOGISIM_NET_230;
   wire s_LOGISIM_NET_231;
   wire s_LOGISIM_NET_232;
   wire s_LOGISIM_NET_233;
   wire s_LOGISIM_NET_234;
   wire s_LOGISIM_NET_235;
   wire s_LOGISIM_NET_236;
   wire s_LOGISIM_NET_237;
   wire s_LOGISIM_NET_238;
   wire s_LOGISIM_NET_239;
   wire s_LOGISIM_NET_24;
   wire s_LOGISIM_NET_240;
   wire s_LOGISIM_NET_241;
   wire s_LOGISIM_NET_242;
   wire s_LOGISIM_NET_243;
   wire s_LOGISIM_NET_244;
   wire s_LOGISIM_NET_245;
   wire s_LOGISIM_NET_246;
   wire s_LOGISIM_NET_247;
   wire s_LOGISIM_NET_248;
   wire s_LOGISIM_NET_249;
   wire s_LOGISIM_NET_25;
   wire s_LOGISIM_NET_250;
   wire s_LOGISIM_NET_251;
   wire s_LOGISIM_NET_252;
   wire s_LOGISIM_NET_253;
   wire s_LOGISIM_NET_254;
   wire s_LOGISIM_NET_255;
   wire s_LOGISIM_NET_256;
   wire s_LOGISIM_NET_257;
   wire s_LOGISIM_NET_258;
   wire s_LOGISIM_NET_259;
   wire s_LOGISIM_NET_26;
   wire s_LOGISIM_NET_260;
   wire s_LOGISIM_NET_261;
   wire s_LOGISIM_NET_262;
   wire s_LOGISIM_NET_263;
   wire s_LOGISIM_NET_264;
   wire s_LOGISIM_NET_265;
   wire s_LOGISIM_NET_266;
   wire s_LOGISIM_NET_267;
   wire s_LOGISIM_NET_27;
   wire s_LOGISIM_NET_28;
   wire s_LOGISIM_NET_29;
   wire s_LOGISIM_NET_3;
   wire s_LOGISIM_NET_30;
   wire s_LOGISIM_NET_31;
   wire s_LOGISIM_NET_32;
   wire s_LOGISIM_NET_33;
   wire s_LOGISIM_NET_34;
   wire s_LOGISIM_NET_35;
   wire s_LOGISIM_NET_36;
   wire s_LOGISIM_NET_37;
   wire s_LOGISIM_NET_38;
   wire s_LOGISIM_NET_39;
   wire s_LOGISIM_NET_4;
   wire s_LOGISIM_NET_40;
   wire s_LOGISIM_NET_41;
   wire s_LOGISIM_NET_42;
   wire s_LOGISIM_NET_43;
   wire s_LOGISIM_NET_44;
   wire s_LOGISIM_NET_45;
   wire s_LOGISIM_NET_46;
   wire s_LOGISIM_NET_47;
   wire s_LOGISIM_NET_48;
   wire s_LOGISIM_NET_49;
   wire s_LOGISIM_NET_5;
   wire s_LOGISIM_NET_50;
   wire s_LOGISIM_NET_51;
   wire s_LOGISIM_NET_52;
   wire s_LOGISIM_NET_53;
   wire s_LOGISIM_NET_54;
   wire s_LOGISIM_NET_55;
   wire s_LOGISIM_NET_56;
   wire s_LOGISIM_NET_57;
   wire s_LOGISIM_NET_58;
   wire s_LOGISIM_NET_59;
   wire s_LOGISIM_NET_6;
   wire s_LOGISIM_NET_60;
   wire s_LOGISIM_NET_61;
   wire s_LOGISIM_NET_62;
   wire s_LOGISIM_NET_63;
   wire s_LOGISIM_NET_64;
   wire s_LOGISIM_NET_65;
   wire s_LOGISIM_NET_66;
   wire s_LOGISIM_NET_67;
   wire s_LOGISIM_NET_68;
   wire s_LOGISIM_NET_69;
   wire s_LOGISIM_NET_7;
   wire s_LOGISIM_NET_70;
   wire s_LOGISIM_NET_71;
   wire s_LOGISIM_NET_72;
   wire s_LOGISIM_NET_73;
   wire s_LOGISIM_NET_74;
   wire s_LOGISIM_NET_75;
   wire s_LOGISIM_NET_76;
   wire s_LOGISIM_NET_77;
   wire s_LOGISIM_NET_78;
   wire s_LOGISIM_NET_79;
   wire s_LOGISIM_NET_8;
   wire s_LOGISIM_NET_80;
   wire s_LOGISIM_NET_81;
   wire s_LOGISIM_NET_82;
   wire s_LOGISIM_NET_83;
   wire s_LOGISIM_NET_84;
   wire s_LOGISIM_NET_85;
   wire s_LOGISIM_NET_86;
   wire s_LOGISIM_NET_87;
   wire s_LOGISIM_NET_88;
   wire s_LOGISIM_NET_89;
   wire s_LOGISIM_NET_9;
   wire s_LOGISIM_NET_90;
   wire s_LOGISIM_NET_91;
   wire s_LOGISIM_NET_92;
   wire s_LOGISIM_NET_93;
   wire s_LOGISIM_NET_94;
   wire s_LOGISIM_NET_95;
   wire s_LOGISIM_NET_96;
   wire s_LOGISIM_NET_97;
   wire s_LOGISIM_NET_98;
   wire s_LOGISIM_NET_99;


   /***************************************************************************
    ** Here all input connections are defined                                **
    ***************************************************************************/
   assign s_LOGISIM_NET_35                   = F30;
   assign s_LOGISIM_NET_14                   = OP5;
   assign s_LOGISIM_NET_29                   = F25;
   assign s_LOGISIM_NET_1                    = OP3;
   assign s_LOGISIM_NET_7                    = OP2;
   assign s_LOGISIM_NET_2                    = OP6;
   assign s_LOGISIM_NET_18                   = OP4;
   assign s_LOGISIM_NET_12                   = F12;
   assign s_LOGISIM_NET_13                   = F14;
   assign s_LOGISIM_NET_28                   = F13;

   /***************************************************************************
    ** Here all output connections are defined                               **
    ***************************************************************************/
   assign half                               = s_LOGISIM_NET_251;
   assign S_Type                             = s_LOGISIM_NET_88;
   assign JAL                                = s_LOGISIM_NET_266;
   assign JALR                               = s_LOGISIM_NET_113;
   assign ALU_SRC                            = s_LOGISIM_NET_143;
   assign BEQ                                = s_LOGISIM_NET_137;
   assign ecall                              = s_LOGISIM_NET_260;
   assign MemWrite                           = s_LOGISIM_NET_122;
   assign BNE                                = s_LOGISIM_NET_226;
   assign CSR                                = s_LOGISIM_NET_223;
   assign RegWrite                           = s_LOGISIM_NET_250;
   assign MemToReg                           = s_LOGISIM_NET_198;

   /***************************************************************************
    ** Here all normal components are defined                                **
    ***************************************************************************/
   NOT_GATE      GATE_1 (.Input_1(s_LOGISIM_NET_1),
                         .Result(s_LOGISIM_NET_78));

   NOT_GATE      GATE_2 (.Input_1(s_LOGISIM_NET_2),
                         .Result(s_LOGISIM_NET_54));

   NOT_GATE      GATE_3 (.Input_1(s_LOGISIM_NET_12),
                         .Result(s_LOGISIM_NET_125));

   NOT_GATE      GATE_4 (.Input_1(s_LOGISIM_NET_28),
                         .Result(s_LOGISIM_NET_77));

   NOT_GATE      GATE_5 (.Input_1(s_LOGISIM_NET_2),
                         .Result(s_LOGISIM_NET_46));

   NOT_GATE      GATE_6 (.Input_1(s_LOGISIM_NET_7),
                         .Result(s_LOGISIM_NET_147));

   NOT_GATE      GATE_7 (.Input_1(s_LOGISIM_NET_1),
                         .Result(s_LOGISIM_NET_59));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_8 (.Input_1(s_LOGISIM_NET_73),
              .Input_2(s_LOGISIM_NET_78),
              .Input_3(s_LOGISIM_NET_18),
              .Input_4(s_LOGISIM_NET_14),
              .Input_5(s_LOGISIM_NET_2),
              .Input_6(s_LOGISIM_NET_28),
              .Input_7(s_LOGISIM_NET_13),
              .Result(s_LOGISIM_NET_221));

   NOT_GATE      GATE_9 (.Input_1(s_LOGISIM_NET_2),
                         .Result(s_LOGISIM_NET_92));

   NOT_GATE      GATE_10 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_216));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_11 (.Input_1(s_LOGISIM_NET_217),
               .Input_10(s_LOGISIM_NET_96),
               .Input_2(s_LOGISIM_NET_149),
               .Input_3(s_LOGISIM_NET_13),
               .Input_4(s_LOGISIM_NET_77),
               .Input_5(s_LOGISIM_NET_180),
               .Input_6(s_LOGISIM_NET_33),
               .Input_7(s_LOGISIM_NET_14),
               .Input_8(s_LOGISIM_NET_18),
               .Input_9(s_LOGISIM_NET_85),
               .Result(s_LOGISIM_NET_58));

   NOT_GATE      GATE_12 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_175));

   NOT_GATE      GATE_13 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_254));

   NOT_GATE      GATE_14 (.Input_1(s_LOGISIM_NET_28),
                          .Result(s_LOGISIM_NET_70));

   NOT_GATE      GATE_15 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_32));

   NOT_GATE      GATE_16 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_261));

   NOT_GATE      GATE_17 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_220));

   NOT_GATE      GATE_18 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_44));

   OR_GATE_20_INPUTS #(.BubblesMask(0))
      GATE_19 (.Input_1(s_LOGISIM_NET_25),
               .Input_10(s_LOGISIM_NET_57),
               .Input_11(s_LOGISIM_NET_207),
               .Input_12(s_LOGISIM_NET_138),
               .Input_13(s_LOGISIM_NET_26),
               .Input_14(s_LOGISIM_NET_82),
               .Input_15(s_LOGISIM_NET_121),
               .Input_16(s_LOGISIM_NET_160),
               .Input_17(s_LOGISIM_NET_190),
               .Input_18(s_LOGISIM_NET_177),
               .Input_19(s_LOGISIM_NET_58),
               .Input_2(s_LOGISIM_NET_60),
               .Input_20(s_LOGISIM_NET_40),
               .Input_3(s_LOGISIM_NET_97),
               .Input_4(s_LOGISIM_NET_168),
               .Input_5(s_LOGISIM_NET_155),
               .Input_6(s_LOGISIM_NET_134),
               .Input_7(s_LOGISIM_NET_206),
               .Input_8(s_LOGISIM_NET_6),
               .Input_9(s_LOGISIM_NET_239),
               .Result(s_LOGISIM_NET_250));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_20 (.Input_1(s_LOGISIM_NET_13),
               .Input_2(s_LOGISIM_NET_28),
               .Input_3(s_LOGISIM_NET_12),
               .Input_4(s_LOGISIM_NET_262),
               .Input_5(s_LOGISIM_NET_232),
               .Input_6(s_LOGISIM_NET_18),
               .Input_7(s_LOGISIM_NET_144),
               .Input_8(s_LOGISIM_NET_81),
               .Result(s_LOGISIM_NET_6));

   NOT_GATE      GATE_21 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_163));

   NOT_GATE      GATE_22 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_124));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_23 (.Input_1(s_LOGISIM_NET_76),
               .Input_2(s_LOGISIM_NET_233),
               .Input_3(s_LOGISIM_NET_18),
               .Input_4(s_LOGISIM_NET_14),
               .Input_5(s_LOGISIM_NET_2),
               .Input_6(s_LOGISIM_NET_28),
               .Input_7(s_LOGISIM_NET_13),
               .Result(s_LOGISIM_NET_223));

   NOT_GATE      GATE_24 (.Input_1(s_LOGISIM_NET_29),
                          .Result(s_LOGISIM_NET_72));

   NOT_GATE      GATE_25 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_262));

   NOT_GATE      GATE_26 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_68));

   NOT_GATE      GATE_27 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_237));

   NOT_GATE      GATE_28 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_67));

   NOT_GATE      GATE_29 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_95));

   NOT_GATE      GATE_30 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_231));

   NOT_GATE      GATE_31 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_214));

   NOT_GATE      GATE_32 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_83));

   NOT_GATE      GATE_33 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_162));

   NOT_GATE      GATE_34 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_108));

   NOT_GATE      GATE_35 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_263));

   NOT_GATE      GATE_36 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_80));

   NOT_GATE      GATE_37 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_90));

   NOT_GATE      GATE_38 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_94));

   NOT_GATE      GATE_39 (.Input_1(s_LOGISIM_NET_28),
                          .Result(s_LOGISIM_NET_188));

   NOT_GATE      GATE_40 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_64));

   NOT_GATE      GATE_41 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_116));

   NOT_GATE      GATE_42 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_265));

   NOT_GATE      GATE_43 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_185));

   NOT_GATE      GATE_44 (.Input_1(s_LOGISIM_NET_28),
                          .Result(s_LOGISIM_NET_103));

   NOT_GATE      GATE_45 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_228));

   NOT_GATE      GATE_46 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_115));

   NOT_GATE      GATE_47 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_167));

   NOT_GATE      GATE_48 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_106));

   NOT_GATE      GATE_49 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_259));

   NOT_GATE      GATE_50 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_76));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_51 (.Input_1(s_LOGISIM_NET_7),
               .Input_2(s_LOGISIM_NET_131),
               .Input_3(s_LOGISIM_NET_248),
               .Input_4(s_LOGISIM_NET_14),
               .Input_5(s_LOGISIM_NET_2),
               .Input_6(s_LOGISIM_NET_169),
               .Input_7(s_LOGISIM_NET_109),
               .Input_8(s_LOGISIM_NET_20),
               .Result(s_LOGISIM_NET_113));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_52 (.Input_1(s_LOGISIM_NET_7),
               .Input_2(s_LOGISIM_NET_59),
               .Input_3(s_LOGISIM_NET_211),
               .Input_4(s_LOGISIM_NET_14),
               .Input_5(s_LOGISIM_NET_2),
               .Input_6(s_LOGISIM_NET_62),
               .Input_7(s_LOGISIM_NET_103),
               .Input_8(s_LOGISIM_NET_219),
               .Result(s_LOGISIM_NET_230));

   NOT_GATE      GATE_53 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_37));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_54 (.Input_1(s_LOGISIM_NET_32),
               .Input_10(s_LOGISIM_NET_167),
               .Input_2(s_LOGISIM_NET_183),
               .Input_3(s_LOGISIM_NET_13),
               .Input_4(s_LOGISIM_NET_243),
               .Input_5(s_LOGISIM_NET_12),
               .Input_6(s_LOGISIM_NET_45),
               .Input_7(s_LOGISIM_NET_153),
               .Input_8(s_LOGISIM_NET_18),
               .Input_9(s_LOGISIM_NET_228),
               .Result(s_LOGISIM_NET_26));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_55 (.Input_1(s_LOGISIM_NET_95),
               .Input_2(s_LOGISIM_NET_255),
               .Input_3(s_LOGISIM_NET_158),
               .Input_4(s_LOGISIM_NET_192),
               .Input_5(s_LOGISIM_NET_52),
               .Input_6(s_LOGISIM_NET_18),
               .Input_7(s_LOGISIM_NET_19),
               .Input_8(s_LOGISIM_NET_178),
               .Result(s_LOGISIM_NET_206));

   NOT_GATE      GATE_56 (.Input_1(s_LOGISIM_NET_29),
                          .Result(s_LOGISIM_NET_174));

   NOT_GATE      GATE_57 (.Input_1(s_LOGISIM_NET_29),
                          .Result(s_LOGISIM_NET_149));

   NOT_GATE      GATE_58 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_128));

   NOT_GATE      GATE_59 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_87));

   NOT_GATE      GATE_60 (.Input_1(s_LOGISIM_NET_28),
                          .Result(s_LOGISIM_NET_9));

   NOT_GATE      GATE_61 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_107));

   NOT_GATE      GATE_62 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_55));

   NOT_GATE      GATE_63 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_187));

   NOT_GATE      GATE_64 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_53));

   NOT_GATE      GATE_65 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_56));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_66 (.Input_1(s_LOGISIM_NET_35),
               .Input_10(s_LOGISIM_NET_94),
               .Input_2(s_LOGISIM_NET_174),
               .Input_3(s_LOGISIM_NET_235),
               .Input_4(s_LOGISIM_NET_79),
               .Input_5(s_LOGISIM_NET_179),
               .Input_6(s_LOGISIM_NET_31),
               .Input_7(s_LOGISIM_NET_14),
               .Input_8(s_LOGISIM_NET_18),
               .Input_9(s_LOGISIM_NET_87),
               .Result(s_LOGISIM_NET_60));

   NOT_GATE      GATE_67 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_3));

   NOT_GATE      GATE_68 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_197));

   NOT_GATE      GATE_69 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_140));

   NOT_GATE      GATE_70 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_10));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_71 (.Input_1(s_LOGISIM_NET_80),
               .Input_10(s_LOGISIM_NET_0),
               .Input_2(s_LOGISIM_NET_120),
               .Input_3(s_LOGISIM_NET_39),
               .Input_4(s_LOGISIM_NET_188),
               .Input_5(s_LOGISIM_NET_236),
               .Input_6(s_LOGISIM_NET_92),
               .Input_7(s_LOGISIM_NET_14),
               .Input_8(s_LOGISIM_NET_18),
               .Input_9(s_LOGISIM_NET_196),
               .Result(s_LOGISIM_NET_25));

   NOT_GATE      GATE_72 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_179));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_73 (.Input_1(s_LOGISIM_NET_162),
               .Input_2(s_LOGISIM_NET_28),
               .Input_3(s_LOGISIM_NET_125),
               .Input_4(s_LOGISIM_NET_164),
               .Input_5(s_LOGISIM_NET_5),
               .Input_6(s_LOGISIM_NET_140),
               .Input_7(s_LOGISIM_NET_141),
               .Input_8(s_LOGISIM_NET_150),
               .Result(s_LOGISIM_NET_121));

   NOT_GATE      GATE_74 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_233));

   NOT_GATE      GATE_75 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_62));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_76 (.Input_1(s_LOGISIM_NET_215),
               .Input_2(s_LOGISIM_NET_67),
               .Input_3(s_LOGISIM_NET_18),
               .Input_4(s_LOGISIM_NET_98),
               .Input_5(s_LOGISIM_NET_24),
               .Input_6(s_LOGISIM_NET_28),
               .Input_7(s_LOGISIM_NET_13),
               .Result(s_LOGISIM_NET_159));

   NOT_GATE      GATE_77 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_4));

   NOT_GATE      GATE_78 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_219));

   NOT_GATE      GATE_79 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_249));

   NOT_GATE      GATE_80 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_153));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_81 (.Input_1(s_LOGISIM_NET_47),
               .Input_2(s_LOGISIM_NET_234),
               .Input_3(s_LOGISIM_NET_36),
               .Input_4(s_LOGISIM_NET_14),
               .Input_5(s_LOGISIM_NET_2),
               .Input_6(s_LOGISIM_NET_12),
               .Input_7(s_LOGISIM_NET_50),
               .Input_8(s_LOGISIM_NET_53),
               .Result(s_LOGISIM_NET_226));

   NOT_GATE      GATE_82 (.Input_1(s_LOGISIM_NET_35),
                          .Result(s_LOGISIM_NET_182));

   NOT_GATE      GATE_83 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_27));

   NOT_GATE      GATE_84 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_49));

   NOT_GATE      GATE_85 (.Input_1(s_LOGISIM_NET_14),
                          .Result(s_LOGISIM_NET_238));

   NOT_GATE      GATE_86 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_73));

   NOT_GATE      GATE_87 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_112));

   NOT_GATE      GATE_88 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_102));

   NOT_GATE      GATE_89 (.Input_1(s_LOGISIM_NET_28),
                          .Result(s_LOGISIM_NET_170));

   NOT_GATE      GATE_90 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_85));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_91 (.Input_1(s_LOGISIM_NET_135),
               .Input_2(s_LOGISIM_NET_146),
               .Input_3(s_LOGISIM_NET_252),
               .Input_4(s_LOGISIM_NET_14),
               .Input_5(s_LOGISIM_NET_83),
               .Input_6(s_LOGISIM_NET_187),
               .Input_7(s_LOGISIM_NET_28),
               .Input_8(s_LOGISIM_NET_42),
               .Result(s_LOGISIM_NET_122));

   NOT_GATE      GATE_92 (.Input_1(s_LOGISIM_NET_12),
                          .Result(s_LOGISIM_NET_241));

   NOT_GATE      GATE_93 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_203));

   NOT_GATE      GATE_94 (.Input_1(s_LOGISIM_NET_18),
                          .Result(s_LOGISIM_NET_184));

   NOT_GATE      GATE_95 (.Input_1(s_LOGISIM_NET_1),
                          .Result(s_LOGISIM_NET_145));

   NOT_GATE      GATE_96 (.Input_1(s_LOGISIM_NET_7),
                          .Result(s_LOGISIM_NET_178));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_97 (.Input_1(s_LOGISIM_NET_86),
               .Input_2(s_LOGISIM_NET_133),
               .Input_3(s_LOGISIM_NET_254),
               .Input_4(s_LOGISIM_NET_259),
               .Input_5(s_LOGISIM_NET_225),
               .Input_6(s_LOGISIM_NET_12),
               .Input_7(s_LOGISIM_NET_129),
               .Input_8(s_LOGISIM_NET_13),
               .Result(s_LOGISIM_NET_227));

   NOT_GATE      GATE_98 (.Input_1(s_LOGISIM_NET_2),
                          .Result(s_LOGISIM_NET_31));

   NOT_GATE      GATE_99 (.Input_1(s_LOGISIM_NET_13),
                          .Result(s_LOGISIM_NET_191));

   NOT_GATE      GATE_100 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_91));

   NOT_GATE      GATE_101 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_181));

   NOT_GATE      GATE_102 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_81));

   NOT_GATE      GATE_103 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_24));

   NOT_GATE      GATE_104 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_5));

   NOT_GATE      GATE_105 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_98));

   NOT_GATE      GATE_106 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_267));

   NOT_GATE      GATE_107 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_17));

   NOT_GATE      GATE_108 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_20));

   NOT_GATE      GATE_109 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_30));

   NOT_GATE      GATE_110 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_247));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_111 (.Input_1(s_LOGISIM_NET_99),
                .Input_10(s_LOGISIM_NET_68),
                .Input_2(s_LOGISIM_NET_151),
                .Input_3(s_LOGISIM_NET_200),
                .Input_4(s_LOGISIM_NET_9),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_163),
                .Input_7(s_LOGISIM_NET_21),
                .Input_8(s_LOGISIM_NET_18),
                .Input_9(s_LOGISIM_NET_128),
                .Result(s_LOGISIM_NET_138));

   NOT_GATE      GATE_112 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_127));

   AND_GATE_6_INPUTS #(.BubblesMask(0))
      GATE_113 (.Input_1(s_LOGISIM_NET_102),
                .Input_2(s_LOGISIM_NET_106),
                .Input_3(s_LOGISIM_NET_18),
                .Input_4(s_LOGISIM_NET_231),
                .Input_5(s_LOGISIM_NET_185),
                .Input_6(s_LOGISIM_NET_114),
                .Result(s_LOGISIM_NET_157));

   NOT_GATE      GATE_114 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_235));

   NOT_GATE      GATE_115 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_139));

   NOT_GATE      GATE_116 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_256));

   NOT_GATE      GATE_117 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_245));

   NOT_GATE      GATE_118 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_104));

   NOT_GATE      GATE_119 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_61));

   NOT_GATE      GATE_120 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_42));

   NOT_GATE      GATE_121 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_211));

   NOT_GATE      GATE_122 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_22));

   NOT_GATE      GATE_123 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_41));

   NOT_GATE      GATE_124 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_135));

   NOT_GATE      GATE_125 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_240));

   NOT_GATE      GATE_126 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_110));

   NOT_GATE      GATE_127 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_16));

   NOT_GATE      GATE_128 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_21));

   NOT_GATE      GATE_129 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_246));

   NOT_GATE      GATE_130 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_34));

   NOT_GATE      GATE_131 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_218));

   NOT_GATE      GATE_132 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_217));

   NOT_GATE      GATE_133 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_243));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_134 (.Input_1(s_LOGISIM_NET_107),
                .Input_10(s_LOGISIM_NET_49),
                .Input_2(s_LOGISIM_NET_72),
                .Input_3(s_LOGISIM_NET_75),
                .Input_4(s_LOGISIM_NET_28),
                .Input_5(s_LOGISIM_NET_241),
                .Input_6(s_LOGISIM_NET_117),
                .Input_7(s_LOGISIM_NET_14),
                .Input_8(s_LOGISIM_NET_18),
                .Input_9(s_LOGISIM_NET_210),
                .Result(s_LOGISIM_NET_155));

   NOT_GATE      GATE_135 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_212));

   NOT_GATE      GATE_136 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_215));

   NOT_GATE      GATE_137 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_45));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_138 (.Input_1(s_LOGISIM_NET_93),
                .Input_10(s_LOGISIM_NET_208),
                .Input_2(s_LOGISIM_NET_8),
                .Input_3(s_LOGISIM_NET_13),
                .Input_4(s_LOGISIM_NET_28),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_264),
                .Input_7(s_LOGISIM_NET_14),
                .Input_8(s_LOGISIM_NET_18),
                .Input_9(s_LOGISIM_NET_136),
                .Result(s_LOGISIM_NET_97));

   NOT_GATE      GATE_139 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_176));

   NOT_GATE      GATE_140 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_33));

   NOT_GATE      GATE_141 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_196));

   NOT_GATE      GATE_142 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_100));

   NOT_GATE      GATE_143 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_253));

   NOT_GATE      GATE_144 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_65));

   NOT_GATE      GATE_145 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_126));

   NOT_GATE      GATE_146 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_166));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_147 (.Input_1(s_LOGISIM_NET_69),
                .Input_2(s_LOGISIM_NET_249),
                .Input_3(s_LOGISIM_NET_124),
                .Input_4(s_LOGISIM_NET_165),
                .Input_5(s_LOGISIM_NET_4),
                .Input_6(s_LOGISIM_NET_12),
                .Input_7(s_LOGISIM_NET_139),
                .Input_8(s_LOGISIM_NET_13),
                .Result(s_LOGISIM_NET_251));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_148 (.Input_1(s_LOGISIM_NET_224),
                .Input_10(s_LOGISIM_NET_44),
                .Input_2(s_LOGISIM_NET_126),
                .Input_3(s_LOGISIM_NET_104),
                .Input_4(s_LOGISIM_NET_28),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_229),
                .Input_7(s_LOGISIM_NET_14),
                .Input_8(s_LOGISIM_NET_18),
                .Input_9(s_LOGISIM_NET_37),
                .Result(s_LOGISIM_NET_134));

   NOT_GATE      GATE_149 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_136));

   NOT_GATE      GATE_150 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_169));

   NOT_GATE      GATE_151 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_258));

   NOT_GATE      GATE_152 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_0));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_153 (.Input_1(s_LOGISIM_NET_41),
                .Input_2(s_LOGISIM_NET_216),
                .Input_3(s_LOGISIM_NET_55),
                .Input_4(s_LOGISIM_NET_48),
                .Input_5(s_LOGISIM_NET_11),
                .Input_6(s_LOGISIM_NET_12),
                .Input_7(s_LOGISIM_NET_15),
                .Input_8(s_LOGISIM_NET_13),
                .Result(s_LOGISIM_NET_101));

   NOT_GATE      GATE_154 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_161));

   NOT_GATE      GATE_155 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_141));

   NOT_GATE      GATE_156 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_86));

   NOT_GATE      GATE_157 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_209));

   NOT_GATE      GATE_158 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_164));

   NOT_GATE      GATE_159 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_119));

   NOT_GATE      GATE_160 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_165));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_161 (.Input_1(s_LOGISIM_NET_152),
                .Input_2(s_LOGISIM_NET_161),
                .Input_3(s_LOGISIM_NET_10),
                .Input_4(s_LOGISIM_NET_14),
                .Input_5(s_LOGISIM_NET_2),
                .Input_6(s_LOGISIM_NET_199),
                .Input_7(s_LOGISIM_NET_132),
                .Input_8(s_LOGISIM_NET_64),
                .Result(s_LOGISIM_NET_137));

   NOT_GATE      GATE_162 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_204));

   NOT_GATE      GATE_163 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_213));

   NOT_GATE      GATE_164 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_109));

   NOT_GATE      GATE_165 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_74));

   NOT_GATE      GATE_166 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_151));

   NOT_GATE      GATE_167 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_50));

   NOT_GATE      GATE_168 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_193));

   NOT_GATE      GATE_169 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_148));

   NOT_GATE      GATE_170 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_146));

   NOT_GATE      GATE_171 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_63));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_172 (.Input_1(s_LOGISIM_NET_13),
                .Input_2(s_LOGISIM_NET_213),
                .Input_3(s_LOGISIM_NET_12),
                .Input_4(s_LOGISIM_NET_267),
                .Input_5(s_LOGISIM_NET_247),
                .Input_6(s_LOGISIM_NET_176),
                .Input_7(s_LOGISIM_NET_203),
                .Input_8(s_LOGISIM_NET_127),
                .Result(s_LOGISIM_NET_40));

   NOT_GATE      GATE_173 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_15));

   NOT_GATE      GATE_174 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_19));

   NOT_GATE      GATE_175 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_180));

   NOT_GATE      GATE_176 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_48));

   NOT_GATE      GATE_177 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_257));

   OR_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_178 (.Input_1(s_LOGISIM_NET_123),
                .Input_2(s_LOGISIM_NET_101),
                .Input_3(s_LOGISIM_NET_157),
                .Input_4(s_LOGISIM_NET_118),
                .Input_5(s_LOGISIM_NET_51),
                .Input_6(s_LOGISIM_NET_159),
                .Input_7(s_LOGISIM_NET_221),
                .Input_8(s_LOGISIM_NET_230),
                .Result(s_LOGISIM_NET_143));

   NOT_GATE      GATE_179 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_225));

   NOT_GATE      GATE_180 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_200));

   NOT_GATE      GATE_181 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_234));

   NOT_GATE      GATE_182 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_120));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_183 (.Input_1(s_LOGISIM_NET_209),
                .Input_2(s_LOGISIM_NET_212),
                .Input_3(s_LOGISIM_NET_66),
                .Input_4(s_LOGISIM_NET_2),
                .Input_5(s_LOGISIM_NET_14),
                .Input_6(s_LOGISIM_NET_22),
                .Input_7(s_LOGISIM_NET_201),
                .Input_8(s_LOGISIM_NET_7),
                .Result(s_LOGISIM_NET_190));

   NOT_GATE      GATE_184 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_232));

   NOT_GATE      GATE_185 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_99));

   NOT_GATE      GATE_186 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_186));

   NOT_GATE      GATE_187 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_75));

   NOT_GATE      GATE_188 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_96));

   NOT_GATE      GATE_189 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_39));

   NOT_GATE      GATE_190 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_158));

   NOT_GATE      GATE_191 (.Input_1(s_LOGISIM_NET_13),
                           .Result(s_LOGISIM_NET_23));

   NOT_GATE      GATE_192 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_194));

   NOT_GATE      GATE_193 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_142));

   NOT_GATE      GATE_194 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_131));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_195 (.Input_1(s_LOGISIM_NET_35),
                .Input_10(s_LOGISIM_NET_147),
                .Input_2(s_LOGISIM_NET_105),
                .Input_3(s_LOGISIM_NET_13),
                .Input_4(s_LOGISIM_NET_70),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_218),
                .Input_7(s_LOGISIM_NET_115),
                .Input_8(s_LOGISIM_NET_18),
                .Input_9(s_LOGISIM_NET_84),
                .Result(s_LOGISIM_NET_82));

   NOT_GATE      GATE_196 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_242));

   NOT_GATE      GATE_197 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_173));

   NOT_GATE      GATE_198 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_236));

   NOT_GATE      GATE_199 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_52));

   NOT_GATE      GATE_200 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_152));

   NOT_GATE      GATE_201 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_133));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_202 (.Input_1(s_LOGISIM_NET_13),
                .Input_2(s_LOGISIM_NET_119),
                .Input_3(s_LOGISIM_NET_253),
                .Input_4(s_LOGISIM_NET_257),
                .Input_5(s_LOGISIM_NET_222),
                .Input_6(s_LOGISIM_NET_18),
                .Input_7(s_LOGISIM_NET_116),
                .Input_8(s_LOGISIM_NET_43),
                .Result(s_LOGISIM_NET_57));

   NOT_GATE      GATE_203 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_150));

   NOT_GATE      GATE_204 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_93));

   NOT_GATE      GATE_205 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_84));

   NOT_GATE      GATE_206 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_210));

   NOT_GATE      GATE_207 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_47));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_208 (.Input_1(s_LOGISIM_NET_148),
                .Input_10(s_LOGISIM_NET_3),
                .Input_2(s_LOGISIM_NET_34),
                .Input_3(s_LOGISIM_NET_90),
                .Input_4(s_LOGISIM_NET_244),
                .Input_5(s_LOGISIM_NET_12),
                .Input_6(s_LOGISIM_NET_46),
                .Input_7(s_LOGISIM_NET_14),
                .Input_8(s_LOGISIM_NET_18),
                .Input_9(s_LOGISIM_NET_195),
                .Result(s_LOGISIM_NET_177));

   NOT_GATE      GATE_209 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_105));

   NOT_GATE      GATE_210 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_208));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_211 (.Input_1(s_LOGISIM_NET_111),
                .Input_2(s_LOGISIM_NET_16),
                .Input_3(s_LOGISIM_NET_171),
                .Input_4(s_LOGISIM_NET_205),
                .Input_5(s_LOGISIM_NET_71),
                .Input_6(s_LOGISIM_NET_186),
                .Input_7(s_LOGISIM_NET_28),
                .Input_8(s_LOGISIM_NET_191),
                .Result(s_LOGISIM_NET_130));

   NOT_GATE      GATE_212 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_156));

   NOT_GATE      GATE_213 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_252));

   NOT_GATE      GATE_214 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_154));

   NOT_GATE      GATE_215 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_38));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_216 (.Input_1(s_LOGISIM_NET_100),
                .Input_2(s_LOGISIM_NET_108),
                .Input_3(s_LOGISIM_NET_240),
                .Input_4(s_LOGISIM_NET_14),
                .Input_5(s_LOGISIM_NET_30),
                .Input_6(s_LOGISIM_NET_142),
                .Input_7(s_LOGISIM_NET_28),
                .Input_8(s_LOGISIM_NET_245),
                .Result(s_LOGISIM_NET_88));

   NOT_GATE      GATE_217 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_132));

   NOT_GATE      GATE_218 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_255));

   AND_GATE_10_INPUTS #(.BubblesMask(0))
      GATE_219 (.Input_1(s_LOGISIM_NET_181),
                .Input_10(s_LOGISIM_NET_166),
                .Input_2(s_LOGISIM_NET_89),
                .Input_3(s_LOGISIM_NET_13),
                .Input_4(s_LOGISIM_NET_28),
                .Input_5(s_LOGISIM_NET_263),
                .Input_6(s_LOGISIM_NET_214),
                .Input_7(s_LOGISIM_NET_14),
                .Input_8(s_LOGISIM_NET_18),
                .Input_9(s_LOGISIM_NET_91),
                .Result(s_LOGISIM_NET_168));

   NOT_GATE      GATE_220 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_264));

   NOT_GATE      GATE_221 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_205));

   NOT_GATE      GATE_222 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_183));

   NOT_GATE      GATE_223 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_43));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_224 (.Input_1(s_LOGISIM_NET_2),
                .Input_2(s_LOGISIM_NET_14),
                .Input_3(s_LOGISIM_NET_184),
                .Input_4(s_LOGISIM_NET_1),
                .Input_5(s_LOGISIM_NET_7),
                .Result(s_LOGISIM_NET_160));

   NOT_GATE      GATE_225 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_89));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_226 (.Input_1(s_LOGISIM_NET_61),
                .Input_2(s_LOGISIM_NET_202),
                .Input_3(s_LOGISIM_NET_17),
                .Input_4(s_LOGISIM_NET_256),
                .Input_5(s_LOGISIM_NET_173),
                .Input_6(s_LOGISIM_NET_28),
                .Input_7(s_LOGISIM_NET_23),
                .Result(s_LOGISIM_NET_123));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_227 (.Input_1(s_LOGISIM_NET_27),
                .Input_2(s_LOGISIM_NET_28),
                .Input_3(s_LOGISIM_NET_261),
                .Input_4(s_LOGISIM_NET_265),
                .Input_5(s_LOGISIM_NET_238),
                .Input_6(s_LOGISIM_NET_18),
                .Input_7(s_LOGISIM_NET_175),
                .Input_8(s_LOGISIM_NET_110),
                .Result(s_LOGISIM_NET_207));

   NOT_GATE      GATE_228 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_248));

   NOT_GATE      GATE_229 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_244));

   NOT_GATE      GATE_230 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_69));

   NOT_GATE      GATE_231 (.Input_1(s_LOGISIM_NET_35),
                           .Result(s_LOGISIM_NET_224));

   NOT_GATE      GATE_232 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_117));

   NOT_GATE      GATE_233 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_36));

   NOT_GATE      GATE_234 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_201));

   NOT_GATE      GATE_235 (.Input_1(s_LOGISIM_NET_14),
                           .Result(s_LOGISIM_NET_222));

   NOT_GATE      GATE_236 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_111));

   NOT_GATE      GATE_237 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_79));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_238 (.Input_1(s_LOGISIM_NET_112),
                .Input_2(s_LOGISIM_NET_154),
                .Input_3(s_LOGISIM_NET_18),
                .Input_4(s_LOGISIM_NET_14),
                .Input_5(s_LOGISIM_NET_2),
                .Input_6(s_LOGISIM_NET_197),
                .Input_7(s_LOGISIM_NET_63),
                .Input_8(s_LOGISIM_NET_204),
                .Result(s_LOGISIM_NET_260));

   OR_GATE #(.BubblesMask(0))
      GATE_239 (.Input_1(s_LOGISIM_NET_130),
                .Input_2(s_LOGISIM_NET_227),
                .Result(s_LOGISIM_NET_198));

   NOT_GATE      GATE_240 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_229));

   NOT_GATE      GATE_241 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_11));

   AND_GATE_7_INPUTS #(.BubblesMask(0))
      GATE_242 (.Input_1(s_LOGISIM_NET_74),
                .Input_2(s_LOGISIM_NET_145),
                .Input_3(s_LOGISIM_NET_18),
                .Input_4(s_LOGISIM_NET_220),
                .Input_5(s_LOGISIM_NET_38),
                .Input_6(s_LOGISIM_NET_13),
                .Input_7(s_LOGISIM_NET_156),
                .Result(s_LOGISIM_NET_51));

   AND_GATE_5_INPUTS #(.BubblesMask(0))
      GATE_243 (.Input_1(s_LOGISIM_NET_7),
                .Input_2(s_LOGISIM_NET_1),
                .Input_3(s_LOGISIM_NET_258),
                .Input_4(s_LOGISIM_NET_14),
                .Input_5(s_LOGISIM_NET_2),
                .Result(s_LOGISIM_NET_266));

   NOT_GATE      GATE_244 (.Input_1(s_LOGISIM_NET_28),
                           .Result(s_LOGISIM_NET_129));

   NOT_GATE      GATE_245 (.Input_1(s_LOGISIM_NET_7),
                           .Result(s_LOGISIM_NET_189));

   NOT_GATE      GATE_246 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_144));

   NOT_GATE      GATE_247 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_172));

   NOT_GATE      GATE_248 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_114));

   NOT_GATE      GATE_249 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_71));

   NOT_GATE      GATE_250 (.Input_1(s_LOGISIM_NET_18),
                           .Result(s_LOGISIM_NET_171));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_251 (.Input_1(s_LOGISIM_NET_189),
                .Input_2(s_LOGISIM_NET_56),
                .Input_3(s_LOGISIM_NET_18),
                .Input_4(s_LOGISIM_NET_193),
                .Input_5(s_LOGISIM_NET_54),
                .Input_6(s_LOGISIM_NET_170),
                .Input_7(s_LOGISIM_NET_172),
                .Input_8(s_LOGISIM_NET_182),
                .Result(s_LOGISIM_NET_118));

   NOT_GATE      GATE_252 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_199));

   NOT_GATE      GATE_253 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_195));

   AND_GATE_8_INPUTS #(.BubblesMask(0))
      GATE_254 (.Input_1(s_LOGISIM_NET_13),
                .Input_2(s_LOGISIM_NET_28),
                .Input_3(s_LOGISIM_NET_237),
                .Input_4(s_LOGISIM_NET_246),
                .Input_5(s_LOGISIM_NET_194),
                .Input_6(s_LOGISIM_NET_18),
                .Input_7(s_LOGISIM_NET_65),
                .Input_8(s_LOGISIM_NET_242),
                .Result(s_LOGISIM_NET_239));

   NOT_GATE      GATE_255 (.Input_1(s_LOGISIM_NET_1),
                           .Result(s_LOGISIM_NET_202));

   NOT_GATE      GATE_256 (.Input_1(s_LOGISIM_NET_2),
                           .Result(s_LOGISIM_NET_192));

   NOT_GATE      GATE_257 (.Input_1(s_LOGISIM_NET_12),
                           .Result(s_LOGISIM_NET_66));

   NOT_GATE      GATE_258 (.Input_1(s_LOGISIM_NET_29),
                           .Result(s_LOGISIM_NET_8));



endmodule
